module q1(a,b,c,d,e,f);
input a,b,c,d,e;
output f;
wire [0:15] Y;
dec4to16 s0 ({a,b,c,d},e,Y);
assign f=Y[1] | Y[3] | Y[6] | Y[7] | Y[9] | Y[14] | Y[15];
endmodule

module dec4to16(w,e,y);
input [3:0] w;
input e;
output reg [0:15] y;
always @(w,e)
begin 
	if (e==0) y=0;
	else 
		case (w)
		0: y=16'b1000000000000000; 1: y=16'b0100000000000000;
		2: y=16'b0010000000000000; 3: y=16'b0001000000000000;
		4: y=16'b0000100000000000; 5: y=16'b0000010000000000;
		6: y=16'b0000001000000000; 7: y=16'b0000000100000000;
		8: y=16'b0000000010000000; 9: y=16'b0000000001000000;
		10: y=16'b0000000000100000; 11: y=16'b0000000000010000;
		12: y=16'b0000000000001000; 13: y=16'b0000000000000100;
		14: y=16'b0000000000000010; 15: y=16'b0000000000000001;
		endcase
end
endmodule
